`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/07/2020 10:04:31 PM
// Design Name: 
// Module Name: FIFO_v1_0
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module FIFO_v1_0(
        input wire AUDIO_DO,
        input wire clk,
        output wire dataReady,
        output wire [7:0] dataOut
    );
    
    
    
    
    
endmodule
